module tb_top ();
    localparam CLK_PERIOD = 10ns;

    logic clk, n_rst;
    logic [7:0] SSEG_CA, SSEG_AN;
    logic [31:0] writeback;


endmodule
