`timescale 1ns / 1ps
module tb_imm_gen ();
    localparam CLK_PERIOD = 10ns;

    logic clk, n_rst;
    logic [31:0] instr, imm_out;   
endmodule