`timescale 1ns / 1ps
module gpio (
    input logic [15:0] SW, writeback,
    input logic [5:0] BTN,
    output logic [15:0] LED,
    output logic [7:0] SSEG_AN, SSEG_CA 
);

endmodule
